
package hls_long_tail_pkg;
    enum {
        conv_fprop1,
        conv_fprop2,
        conv_fprop3,
        max_pooling_fprop1,
        max_pooling_fprop2,
        fully_connected_fprop
    } hls_enum_t;
    localparam HLS_NUM = 6;
    localparam HLS_CACHE = 0;
    localparam HLS_PARENT = 0;
    localparam [$clog2(HLS_NUM)-1:0] HLS_PARENT_IDX[HLS_PARENT] = {

    };


    //xmem desc
    //alias:input_layer_map_w = input_layer.map_w
    //alias:input_layer_map_h = input_layer.map_h
    //alias:input_layer_map_count = input_layer.map_count
    //alias:input_layer_map = input_layer.map
    //alias:input_layer_kernel_w = input_layer.kernel_w
    //alias:input_layer_kernel_h = input_layer.kernel_h
    //alias:input_layer_kernel_count = input_layer.kernel_count
    //alias:input_layer_kernel = input_layer.kernel
    //alias:input_layer_map_common = input_layer.map_common
    //alias:c1_conv_layer_map_w = c1_conv_layer.map_w
    //alias:c1_conv_layer_map_h = c1_conv_layer.map_h
    //alias:c1_conv_layer_map_count = c1_conv_layer.map_count
    //alias:c1_conv_layer_map = c1_conv_layer.map
    //alias:c1_conv_layer_kernel_w = c1_conv_layer.kernel_w
    //alias:c1_conv_layer_kernel_h = c1_conv_layer.kernel_h
    //alias:c1_conv_layer_kernel_count = c1_conv_layer.kernel_count
    //alias:c1_conv_layer_kernel = c1_conv_layer.kernel
    //alias:c1_conv_layer_map_common = c1_conv_layer.map_common
    //alias:s2_pooling_layer_map_w = s2_pooling_layer.map_w
    //alias:s2_pooling_layer_map_h = s2_pooling_layer.map_h
    //alias:s2_pooling_layer_map_count = s2_pooling_layer.map_count
    //alias:s2_pooling_layer_map = s2_pooling_layer.map
    //alias:s2_pooling_layer_kernel_w = s2_pooling_layer.kernel_w
    //alias:s2_pooling_layer_kernel_h = s2_pooling_layer.kernel_h
    //alias:s2_pooling_layer_kernel_count = s2_pooling_layer.kernel_count
    //alias:s2_pooling_layer_kernel = s2_pooling_layer.kernel
    //alias:s2_pooling_layer_map_common = s2_pooling_layer.map_common
    //alias:c3_conv_layer_map_w = c3_conv_layer.map_w
    //alias:c3_conv_layer_map_h = c3_conv_layer.map_h
    //alias:c3_conv_layer_map_count = c3_conv_layer.map_count
    //alias:c3_conv_layer_map = c3_conv_layer.map
    //alias:c3_conv_layer_kernel_w = c3_conv_layer.kernel_w
    //alias:c3_conv_layer_kernel_h = c3_conv_layer.kernel_h
    //alias:c3_conv_layer_kernel_count = c3_conv_layer.kernel_count
    //alias:c3_conv_layer_kernel = c3_conv_layer.kernel
    //alias:c3_conv_layer_map_common = c3_conv_layer.map_common
    //alias:s4_pooling_layer_map_w = s4_pooling_layer.map_w
    //alias:s4_pooling_layer_map_h = s4_pooling_layer.map_h
    //alias:s4_pooling_layer_map_count = s4_pooling_layer.map_count
    //alias:s4_pooling_layer_map = s4_pooling_layer.map
    //alias:s4_pooling_layer_kernel_w = s4_pooling_layer.kernel_w
    //alias:s4_pooling_layer_kernel_h = s4_pooling_layer.kernel_h
    //alias:s4_pooling_layer_kernel_count = s4_pooling_layer.kernel_count
    //alias:s4_pooling_layer_kernel = s4_pooling_layer.kernel
    //alias:s4_pooling_layer_map_common = s4_pooling_layer.map_common
    //alias:c5_conv_layer_map_w = c5_conv_layer.map_w
    //alias:c5_conv_layer_map_h = c5_conv_layer.map_h
    //alias:c5_conv_layer_map_count = c5_conv_layer.map_count
    //alias:c5_conv_layer_map = c5_conv_layer.map
    //alias:c5_conv_layer_kernel_w = c5_conv_layer.kernel_w
    //alias:c5_conv_layer_kernel_h = c5_conv_layer.kernel_h
    //alias:c5_conv_layer_kernel_count = c5_conv_layer.kernel_count
    //alias:c5_conv_layer_kernel = c5_conv_layer.kernel
    //alias:c5_conv_layer_map_common = c5_conv_layer.map_common
    //alias:output_layer_map_w = output_layer.map_w
    //alias:output_layer_map_h = output_layer.map_h
    //alias:output_layer_map_count = output_layer.map_count
    //alias:output_layer_map = output_layer.map
    //alias:output_layer_kernel_w = output_layer.kernel_w
    //alias:output_layer_kernel_h = output_layer.kernel_h
    //alias:output_layer_kernel_count = output_layer.kernel_count
    //alias:output_layer_kernel = output_layer.kernel
    //alias:output_layer_map_common = output_layer.map_common

    //xmem width
    localparam width_in_data                                       = 64;
    localparam width_in_w                                          = 32;
    localparam width_in_h                                          = 32;
    localparam width_kernel                                        = 64;
    localparam width_kernel_w                                      = 32;
    localparam width_kernel_h                                      = 32;
    localparam width_out_data                                      = 64;
    localparam width_out_w                                         = 32;
    localparam width_out_h                                         = 32;
    //struct:localparam width_input_layer                                   = 21953728;
    localparam width_input_layer_map_w                             = 32;
    localparam width_input_layer_map_h                             = 32;
    localparam width_input_layer_map_count                         = 32;
    //struct:localparam width_input_layer_map                               = 131200;
    localparam width_input_layer_kernel_w                          = 32;
    localparam width_input_layer_kernel_h                          = 32;
    localparam width_input_layer_kernel_count                      = 32;
    //struct:localparam width_input_layer_kernel                            = 3200;
    localparam width_input_layer_map_common                        = 64;
    //struct:localparam width_c1_conv_layer                                 = 21953728;
    localparam width_c1_conv_layer_map_w                           = 32;
    localparam width_c1_conv_layer_map_h                           = 32;
    localparam width_c1_conv_layer_map_count                       = 32;
    //struct:localparam width_c1_conv_layer_map                             = 131200;
    localparam width_c1_conv_layer_kernel_w                        = 32;
    localparam width_c1_conv_layer_kernel_h                        = 32;
    localparam width_c1_conv_layer_kernel_count                    = 32;
    //struct:localparam width_c1_conv_layer_kernel                          = 3200;
    localparam width_c1_conv_layer_map_common                      = 64;
    //struct:localparam width_s2_pooling_layer                              = 21953728;
    localparam width_s2_pooling_layer_map_w                        = 32;
    localparam width_s2_pooling_layer_map_h                        = 32;
    localparam width_s2_pooling_layer_map_count                    = 32;
    //struct:localparam width_s2_pooling_layer_map                          = 131200;
    localparam width_s2_pooling_layer_kernel_w                     = 32;
    localparam width_s2_pooling_layer_kernel_h                     = 32;
    localparam width_s2_pooling_layer_kernel_count                 = 32;
    //struct:localparam width_s2_pooling_layer_kernel                       = 3200;
    localparam width_s2_pooling_layer_map_common                   = 64;
    //struct:localparam width_c3_conv_layer                                 = 21953728;
    localparam width_c3_conv_layer_map_w                           = 32;
    localparam width_c3_conv_layer_map_h                           = 32;
    localparam width_c3_conv_layer_map_count                       = 32;
    //struct:localparam width_c3_conv_layer_map                             = 131200;
    localparam width_c3_conv_layer_kernel_w                        = 32;
    localparam width_c3_conv_layer_kernel_h                        = 32;
    localparam width_c3_conv_layer_kernel_count                    = 32;
    //struct:localparam width_c3_conv_layer_kernel                          = 3200;
    localparam width_c3_conv_layer_map_common                      = 64;
    //struct:localparam width_s4_pooling_layer                              = 21953728;
    localparam width_s4_pooling_layer_map_w                        = 32;
    localparam width_s4_pooling_layer_map_h                        = 32;
    localparam width_s4_pooling_layer_map_count                    = 32;
    //struct:localparam width_s4_pooling_layer_map                          = 131200;
    localparam width_s4_pooling_layer_kernel_w                     = 32;
    localparam width_s4_pooling_layer_kernel_h                     = 32;
    localparam width_s4_pooling_layer_kernel_count                 = 32;
    //struct:localparam width_s4_pooling_layer_kernel                       = 3200;
    localparam width_s4_pooling_layer_map_common                   = 64;
    //struct:localparam width_c5_conv_layer                                 = 21953728;
    localparam width_c5_conv_layer_map_w                           = 32;
    localparam width_c5_conv_layer_map_h                           = 32;
    localparam width_c5_conv_layer_map_count                       = 32;
    //struct:localparam width_c5_conv_layer_map                             = 131200;
    localparam width_c5_conv_layer_kernel_w                        = 32;
    localparam width_c5_conv_layer_kernel_h                        = 32;
    localparam width_c5_conv_layer_kernel_count                    = 32;
    //struct:localparam width_c5_conv_layer_kernel                          = 3200;
    localparam width_c5_conv_layer_map_common                      = 64;
    //struct:localparam width_output_layer                                  = 21953728;
    localparam width_output_layer_map_w                            = 32;
    localparam width_output_layer_map_h                            = 32;
    localparam width_output_layer_map_count                        = 32;
    //struct:localparam width_output_layer_map                              = 131200;
    localparam width_output_layer_kernel_w                         = 32;
    localparam width_output_layer_kernel_h                         = 32;
    localparam width_output_layer_kernel_count                     = 32;
    //struct:localparam width_output_layer_kernel                           = 3200;
    localparam width_output_layer_map_common                       = 64;
    localparam width_pconnection                                   = 8;
    localparam width_xxxxx_paddingA                                = 8;
    localparam width_generic_xmem32                                = 32;

    //xmem offset
    localparam offset_in_data                                      = 0;
    localparam offset_in_w                                         = 8192;
    localparam offset_in_h                                         = 8196;
    localparam offset_kernel                                       = 8200;
    localparam offset_kernel_w                                     = 8400;
    localparam offset_kernel_h                                     = 8404;
    localparam offset_out_data                                     = 8408;
    localparam offset_out_w                                        = 16600;
    localparam offset_out_h                                        = 16604;
    //struct:localparam offset_input_layer                                  = 16608;
    localparam offset_input_layer_map_w                            = 16608;
    localparam offset_input_layer_map_h                            = 16612;
    localparam offset_input_layer_map_count                        = 16616;
    //struct:localparam offset_input_layer_map                              = 16620;
    localparam offset_input_layer_kernel_w                         = 1984620;
    localparam offset_input_layer_kernel_h                         = 1984624;
    localparam offset_input_layer_kernel_count                     = 1984628;
    //struct:localparam offset_input_layer_kernel                           = 1984632;
    localparam offset_input_layer_map_common                       = 2752632;
    //struct:localparam offset_c1_conv_layer                                = 2760824;
    localparam offset_c1_conv_layer_map_w                          = 2760824;
    localparam offset_c1_conv_layer_map_h                          = 2760828;
    localparam offset_c1_conv_layer_map_count                      = 2760832;
    //struct:localparam offset_c1_conv_layer_map                            = 2760836;
    localparam offset_c1_conv_layer_kernel_w                       = 4728836;
    localparam offset_c1_conv_layer_kernel_h                       = 4728840;
    localparam offset_c1_conv_layer_kernel_count                   = 4728844;
    //struct:localparam offset_c1_conv_layer_kernel                         = 4728848;
    localparam offset_c1_conv_layer_map_common                     = 5496848;
    //struct:localparam offset_s2_pooling_layer                             = 5505040;
    localparam offset_s2_pooling_layer_map_w                       = 5505040;
    localparam offset_s2_pooling_layer_map_h                       = 5505044;
    localparam offset_s2_pooling_layer_map_count                   = 5505048;
    //struct:localparam offset_s2_pooling_layer_map                         = 5505052;
    localparam offset_s2_pooling_layer_kernel_w                    = 7473052;
    localparam offset_s2_pooling_layer_kernel_h                    = 7473056;
    localparam offset_s2_pooling_layer_kernel_count                = 7473060;
    //struct:localparam offset_s2_pooling_layer_kernel                      = 7473064;
    localparam offset_s2_pooling_layer_map_common                  = 8241064;
    //struct:localparam offset_c3_conv_layer                                = 8249256;
    localparam offset_c3_conv_layer_map_w                          = 8249256;
    localparam offset_c3_conv_layer_map_h                          = 8249260;
    localparam offset_c3_conv_layer_map_count                      = 8249264;
    //struct:localparam offset_c3_conv_layer_map                            = 8249268;
    localparam offset_c3_conv_layer_kernel_w                       = 10217268;
    localparam offset_c3_conv_layer_kernel_h                       = 10217272;
    localparam offset_c3_conv_layer_kernel_count                   = 10217276;
    //struct:localparam offset_c3_conv_layer_kernel                         = 10217280;
    localparam offset_c3_conv_layer_map_common                     = 10985280;
    //struct:localparam offset_s4_pooling_layer                             = 10993472;
    localparam offset_s4_pooling_layer_map_w                       = 10993472;
    localparam offset_s4_pooling_layer_map_h                       = 10993476;
    localparam offset_s4_pooling_layer_map_count                   = 10993480;
    //struct:localparam offset_s4_pooling_layer_map                         = 10993484;
    localparam offset_s4_pooling_layer_kernel_w                    = 12961484;
    localparam offset_s4_pooling_layer_kernel_h                    = 12961488;
    localparam offset_s4_pooling_layer_kernel_count                = 12961492;
    //struct:localparam offset_s4_pooling_layer_kernel                      = 12961496;
    localparam offset_s4_pooling_layer_map_common                  = 13729496;
    //struct:localparam offset_c5_conv_layer                                = 13737688;
    localparam offset_c5_conv_layer_map_w                          = 13737688;
    localparam offset_c5_conv_layer_map_h                          = 13737692;
    localparam offset_c5_conv_layer_map_count                      = 13737696;
    //struct:localparam offset_c5_conv_layer_map                            = 13737700;
    localparam offset_c5_conv_layer_kernel_w                       = 15705700;
    localparam offset_c5_conv_layer_kernel_h                       = 15705704;
    localparam offset_c5_conv_layer_kernel_count                   = 15705708;
    //struct:localparam offset_c5_conv_layer_kernel                         = 15705712;
    localparam offset_c5_conv_layer_map_common                     = 16473712;
    //struct:localparam offset_output_layer                                 = 16481904;
    localparam offset_output_layer_map_w                           = 16481904;
    localparam offset_output_layer_map_h                           = 16481908;
    localparam offset_output_layer_map_count                       = 16481912;
    //struct:localparam offset_output_layer_map                             = 16481916;
    localparam offset_output_layer_kernel_w                        = 18449916;
    localparam offset_output_layer_kernel_h                        = 18449920;
    localparam offset_output_layer_kernel_count                    = 18449924;
    //struct:localparam offset_output_layer_kernel                          = 18449928;
    localparam offset_output_layer_map_common                      = 19217928;
    localparam offset_pconnection                                  = 19226120;
    localparam offset_xxxxx_paddingA                               = 19226216;
    localparam offset_generic_xmem32                               = 0;

    //xmem depth
    localparam depth_in_data                                       = 1024;
    localparam depth_in_w                                          = 1;
    localparam depth_in_h                                          = 1;
    localparam depth_kernel                                        = 25;
    localparam depth_kernel_w                                      = 1;
    localparam depth_kernel_h                                      = 1;
    localparam depth_out_data                                      = 1024;
    localparam depth_out_w                                         = 1;
    localparam depth_out_h                                         = 1;
    //struct:localparam depth_input_layer                                   = 1;
    localparam depth_input_layer_map_w                             = 1;
    localparam depth_input_layer_map_h                             = 1;
    localparam depth_input_layer_map_count                         = 1;
    //struct:localparam depth_input_layer_map                               = 120;
    localparam depth_input_layer_kernel_w                          = 1;
    localparam depth_input_layer_kernel_h                          = 1;
    localparam depth_input_layer_kernel_count                      = 1;
    //struct:localparam depth_input_layer_kernel                            = 1920;
    localparam depth_input_layer_map_common                        = 1024;
    //struct:localparam depth_c1_conv_layer                                 = 1;
    localparam depth_c1_conv_layer_map_w                           = 1;
    localparam depth_c1_conv_layer_map_h                           = 1;
    localparam depth_c1_conv_layer_map_count                       = 1;
    //struct:localparam depth_c1_conv_layer_map                             = 120;
    localparam depth_c1_conv_layer_kernel_w                        = 1;
    localparam depth_c1_conv_layer_kernel_h                        = 1;
    localparam depth_c1_conv_layer_kernel_count                    = 1;
    //struct:localparam depth_c1_conv_layer_kernel                          = 1920;
    localparam depth_c1_conv_layer_map_common                      = 1024;
    //struct:localparam depth_s2_pooling_layer                              = 1;
    localparam depth_s2_pooling_layer_map_w                        = 1;
    localparam depth_s2_pooling_layer_map_h                        = 1;
    localparam depth_s2_pooling_layer_map_count                    = 1;
    //struct:localparam depth_s2_pooling_layer_map                          = 120;
    localparam depth_s2_pooling_layer_kernel_w                     = 1;
    localparam depth_s2_pooling_layer_kernel_h                     = 1;
    localparam depth_s2_pooling_layer_kernel_count                 = 1;
    //struct:localparam depth_s2_pooling_layer_kernel                       = 1920;
    localparam depth_s2_pooling_layer_map_common                   = 1024;
    //struct:localparam depth_c3_conv_layer                                 = 1;
    localparam depth_c3_conv_layer_map_w                           = 1;
    localparam depth_c3_conv_layer_map_h                           = 1;
    localparam depth_c3_conv_layer_map_count                       = 1;
    //struct:localparam depth_c3_conv_layer_map                             = 120;
    localparam depth_c3_conv_layer_kernel_w                        = 1;
    localparam depth_c3_conv_layer_kernel_h                        = 1;
    localparam depth_c3_conv_layer_kernel_count                    = 1;
    //struct:localparam depth_c3_conv_layer_kernel                          = 1920;
    localparam depth_c3_conv_layer_map_common                      = 1024;
    //struct:localparam depth_s4_pooling_layer                              = 1;
    localparam depth_s4_pooling_layer_map_w                        = 1;
    localparam depth_s4_pooling_layer_map_h                        = 1;
    localparam depth_s4_pooling_layer_map_count                    = 1;
    //struct:localparam depth_s4_pooling_layer_map                          = 120;
    localparam depth_s4_pooling_layer_kernel_w                     = 1;
    localparam depth_s4_pooling_layer_kernel_h                     = 1;
    localparam depth_s4_pooling_layer_kernel_count                 = 1;
    //struct:localparam depth_s4_pooling_layer_kernel                       = 1920;
    localparam depth_s4_pooling_layer_map_common                   = 1024;
    //struct:localparam depth_c5_conv_layer                                 = 1;
    localparam depth_c5_conv_layer_map_w                           = 1;
    localparam depth_c5_conv_layer_map_h                           = 1;
    localparam depth_c5_conv_layer_map_count                       = 1;
    //struct:localparam depth_c5_conv_layer_map                             = 120;
    localparam depth_c5_conv_layer_kernel_w                        = 1;
    localparam depth_c5_conv_layer_kernel_h                        = 1;
    localparam depth_c5_conv_layer_kernel_count                    = 1;
    //struct:localparam depth_c5_conv_layer_kernel                          = 1920;
    localparam depth_c5_conv_layer_map_common                      = 1024;
    //struct:localparam depth_output_layer                                  = 1;
    localparam depth_output_layer_map_w                            = 1;
    localparam depth_output_layer_map_h                            = 1;
    localparam depth_output_layer_map_count                        = 1;
    //struct:localparam depth_output_layer_map                              = 120;
    localparam depth_output_layer_kernel_w                         = 1;
    localparam depth_output_layer_kernel_h                         = 1;
    localparam depth_output_layer_kernel_count                     = 1;
    //struct:localparam depth_output_layer_kernel                           = 1920;
    localparam depth_output_layer_map_common                       = 1024;
    localparam depth_pconnection                                   = 96;
    localparam depth_xxxxx_paddingA                                = 1976;
    localparam depth_generic_xmem32                                = 4807048;

endpackage


package hls_long_tail_pkg;
    enum {
        conv_fprop1,
        conv_fprop2,
        conv_fprop3,
        max_pooling_fprop1,
        max_pooling_fprop2,
        fully_connected_fprop
    } hls_enum_t;
    localparam HLS_NUM = 6;
    localparam HLS_CACHE = 0;
    localparam HLS_PARENT = 0;
    localparam [$clog2(HLS_NUM)-1:0] HLS_PARENT_IDX[HLS_PARENT] = {

    };


    //xmem desc
    //alias:input_layer1_map_w = input_layer1.map_w
    //alias:input_layer1_map_h = input_layer1.map_h
    //alias:input_layer1_map_count = input_layer1.map_count
    //alias:input_layer1_kernel_w = input_layer1.kernel_w
    //alias:input_layer1_kernel_h = input_layer1.kernel_h
    //alias:input_layer1_kernel_count = input_layer1.kernel_count
    //alias:c1_conv_layer1_map_w = c1_conv_layer1.map_w
    //alias:c1_conv_layer1_map_h = c1_conv_layer1.map_h
    //alias:c1_conv_layer1_map_count = c1_conv_layer1.map_count
    //alias:c1_conv_layer1_kernel_w = c1_conv_layer1.kernel_w
    //alias:c1_conv_layer1_kernel_h = c1_conv_layer1.kernel_h
    //alias:c1_conv_layer1_kernel_count = c1_conv_layer1.kernel_count
    //alias:s2_pooling_layer1_map_w = s2_pooling_layer1.map_w
    //alias:s2_pooling_layer1_map_h = s2_pooling_layer1.map_h
    //alias:s2_pooling_layer1_map_count = s2_pooling_layer1.map_count
    //alias:s2_pooling_layer1_kernel_w = s2_pooling_layer1.kernel_w
    //alias:s2_pooling_layer1_kernel_h = s2_pooling_layer1.kernel_h
    //alias:s2_pooling_layer1_kernel_count = s2_pooling_layer1.kernel_count
    //alias:c3_conv_layer1_map_w = c3_conv_layer1.map_w
    //alias:c3_conv_layer1_map_h = c3_conv_layer1.map_h
    //alias:c3_conv_layer1_map_count = c3_conv_layer1.map_count
    //alias:c3_conv_layer1_kernel_w = c3_conv_layer1.kernel_w
    //alias:c3_conv_layer1_kernel_h = c3_conv_layer1.kernel_h
    //alias:c3_conv_layer1_kernel_count = c3_conv_layer1.kernel_count
    //alias:s4_pooling_layer1_map_w = s4_pooling_layer1.map_w
    //alias:s4_pooling_layer1_map_h = s4_pooling_layer1.map_h
    //alias:s4_pooling_layer1_map_count = s4_pooling_layer1.map_count
    //alias:s4_pooling_layer1_kernel_w = s4_pooling_layer1.kernel_w
    //alias:s4_pooling_layer1_kernel_h = s4_pooling_layer1.kernel_h
    //alias:s4_pooling_layer1_kernel_count = s4_pooling_layer1.kernel_count
    //alias:c5_conv_layer1_map_w = c5_conv_layer1.map_w
    //alias:c5_conv_layer1_map_h = c5_conv_layer1.map_h
    //alias:c5_conv_layer1_map_count = c5_conv_layer1.map_count
    //alias:c5_conv_layer1_kernel_w = c5_conv_layer1.kernel_w
    //alias:c5_conv_layer1_kernel_h = c5_conv_layer1.kernel_h
    //alias:c5_conv_layer1_kernel_count = c5_conv_layer1.kernel_count
    //alias:output_layer1_map_w = output_layer1.map_w
    //alias:output_layer1_map_h = output_layer1.map_h
    //alias:output_layer1_map_count = output_layer1.map_count
    //alias:output_layer1_kernel_w = output_layer1.kernel_w
    //alias:output_layer1_kernel_h = output_layer1.kernel_h
    //alias:output_layer1_kernel_count = output_layer1.kernel_count
    //alias:input_layer2_data = input_layer2.data
    //alias:input_layer2_error = input_layer2.error
    //alias:input_layer2_b = input_layer2.b
    //alias:input_layer2_db = input_layer2.db
    //alias:input_layer2_W = input_layer2.W
    //alias:input_layer2_dW = input_layer2.dW
    //alias:input_layer2_map_common = input_layer2.map_common
    //alias:c1_conv_layer2_data = c1_conv_layer2.data
    //alias:c1_conv_layer2_error = c1_conv_layer2.error
    //alias:c1_conv_layer2_b = c1_conv_layer2.b
    //alias:c1_conv_layer2_db = c1_conv_layer2.db
    //alias:c1_conv_layer2_W = c1_conv_layer2.W
    //alias:c1_conv_layer2_dW = c1_conv_layer2.dW
    //alias:c1_conv_layer2_map_common = c1_conv_layer2.map_common
    //alias:s2_pooling_layer2_data = s2_pooling_layer2.data
    //alias:s2_pooling_layer2_error = s2_pooling_layer2.error
    //alias:s2_pooling_layer2_b = s2_pooling_layer2.b
    //alias:s2_pooling_layer2_db = s2_pooling_layer2.db
    //alias:s2_pooling_layer2_W = s2_pooling_layer2.W
    //alias:s2_pooling_layer2_dW = s2_pooling_layer2.dW
    //alias:s2_pooling_layer2_map_common = s2_pooling_layer2.map_common
    //alias:c3_conv_layer2_data = c3_conv_layer2.data
    //alias:c3_conv_layer2_error = c3_conv_layer2.error
    //alias:c3_conv_layer2_b = c3_conv_layer2.b
    //alias:c3_conv_layer2_db = c3_conv_layer2.db
    //alias:c3_conv_layer2_W = c3_conv_layer2.W
    //alias:c3_conv_layer2_dW = c3_conv_layer2.dW
    //alias:c3_conv_layer2_map_common = c3_conv_layer2.map_common
    //alias:s4_pooling_layer2_data = s4_pooling_layer2.data
    //alias:s4_pooling_layer2_error = s4_pooling_layer2.error
    //alias:s4_pooling_layer2_b = s4_pooling_layer2.b
    //alias:s4_pooling_layer2_db = s4_pooling_layer2.db
    //alias:s4_pooling_layer2_W = s4_pooling_layer2.W
    //alias:s4_pooling_layer2_dW = s4_pooling_layer2.dW
    //alias:s4_pooling_layer2_map_common = s4_pooling_layer2.map_common
    //alias:c5_conv_layer2_data = c5_conv_layer2.data
    //alias:c5_conv_layer2_error = c5_conv_layer2.error
    //alias:c5_conv_layer2_b = c5_conv_layer2.b
    //alias:c5_conv_layer2_db = c5_conv_layer2.db
    //alias:c5_conv_layer2_W = c5_conv_layer2.W
    //alias:c5_conv_layer2_dW = c5_conv_layer2.dW
    //alias:c5_conv_layer2_map_common = c5_conv_layer2.map_common
    //alias:output_layer2_data = output_layer2.data
    //alias:output_layer2_error = output_layer2.error
    //alias:output_layer2_b = output_layer2.b
    //alias:output_layer2_db = output_layer2.db
    //alias:output_layer2_W = output_layer2.W
    //alias:output_layer2_dW = output_layer2.dW
    //alias:output_layer2_map_common = output_layer2.map_common

    //xmem width
    //struct:localparam width_input_layer1                                  = 192;
    localparam width_input_layer1_map_w                            = 32;
    localparam width_input_layer1_map_h                            = 32;
    localparam width_input_layer1_map_count                        = 32;
    localparam width_input_layer1_kernel_w                         = 32;
    localparam width_input_layer1_kernel_h                         = 32;
    localparam width_input_layer1_kernel_count                     = 32;
    //struct:localparam width_c1_conv_layer1                                = 192;
    localparam width_c1_conv_layer1_map_w                          = 32;
    localparam width_c1_conv_layer1_map_h                          = 32;
    localparam width_c1_conv_layer1_map_count                      = 32;
    localparam width_c1_conv_layer1_kernel_w                       = 32;
    localparam width_c1_conv_layer1_kernel_h                       = 32;
    localparam width_c1_conv_layer1_kernel_count                   = 32;
    //struct:localparam width_s2_pooling_layer1                             = 192;
    localparam width_s2_pooling_layer1_map_w                       = 32;
    localparam width_s2_pooling_layer1_map_h                       = 32;
    localparam width_s2_pooling_layer1_map_count                   = 32;
    localparam width_s2_pooling_layer1_kernel_w                    = 32;
    localparam width_s2_pooling_layer1_kernel_h                    = 32;
    localparam width_s2_pooling_layer1_kernel_count                = 32;
    //struct:localparam width_c3_conv_layer1                                = 192;
    localparam width_c3_conv_layer1_map_w                          = 32;
    localparam width_c3_conv_layer1_map_h                          = 32;
    localparam width_c3_conv_layer1_map_count                      = 32;
    localparam width_c3_conv_layer1_kernel_w                       = 32;
    localparam width_c3_conv_layer1_kernel_h                       = 32;
    localparam width_c3_conv_layer1_kernel_count                   = 32;
    //struct:localparam width_s4_pooling_layer1                             = 192;
    localparam width_s4_pooling_layer1_map_w                       = 32;
    localparam width_s4_pooling_layer1_map_h                       = 32;
    localparam width_s4_pooling_layer1_map_count                   = 32;
    localparam width_s4_pooling_layer1_kernel_w                    = 32;
    localparam width_s4_pooling_layer1_kernel_h                    = 32;
    localparam width_s4_pooling_layer1_kernel_count                = 32;
    //struct:localparam width_c5_conv_layer1                                = 192;
    localparam width_c5_conv_layer1_map_w                          = 32;
    localparam width_c5_conv_layer1_map_h                          = 32;
    localparam width_c5_conv_layer1_map_count                      = 32;
    localparam width_c5_conv_layer1_kernel_w                       = 32;
    localparam width_c5_conv_layer1_kernel_h                       = 32;
    localparam width_c5_conv_layer1_kernel_count                   = 32;
    //struct:localparam width_output_layer1                                 = 192;
    localparam width_output_layer1_map_w                           = 32;
    localparam width_output_layer1_map_h                           = 32;
    localparam width_output_layer1_map_count                       = 32;
    localparam width_output_layer1_kernel_w                        = 32;
    localparam width_output_layer1_kernel_h                        = 32;
    localparam width_output_layer1_kernel_count                    = 32;
    localparam width_xxxxx_paddingA                                = 8;
    //struct:localparam width_input_layer2                                  = 21953536;
    localparam width_input_layer2_data                             = 64;
    localparam width_input_layer2_error                            = 64;
    localparam width_input_layer2_b                                = 64;
    localparam width_input_layer2_db                               = 64;
    localparam width_input_layer2_W                                = 64;
    localparam width_input_layer2_dW                               = 64;
    localparam width_input_layer2_map_common                       = 64;
    //struct:localparam width_c1_conv_layer2                                = 21953536;
    localparam width_c1_conv_layer2_data                           = 64;
    localparam width_c1_conv_layer2_error                          = 64;
    localparam width_c1_conv_layer2_b                              = 64;
    localparam width_c1_conv_layer2_db                             = 64;
    localparam width_c1_conv_layer2_W                              = 64;
    localparam width_c1_conv_layer2_dW                             = 64;
    localparam width_c1_conv_layer2_map_common                     = 64;
    //struct:localparam width_s2_pooling_layer2                             = 21953536;
    localparam width_s2_pooling_layer2_data                        = 64;
    localparam width_s2_pooling_layer2_error                       = 64;
    localparam width_s2_pooling_layer2_b                           = 64;
    localparam width_s2_pooling_layer2_db                          = 64;
    localparam width_s2_pooling_layer2_W                           = 64;
    localparam width_s2_pooling_layer2_dW                          = 64;
    localparam width_s2_pooling_layer2_map_common                  = 64;
    //struct:localparam width_c3_conv_layer2                                = 21953536;
    localparam width_c3_conv_layer2_data                           = 64;
    localparam width_c3_conv_layer2_error                          = 64;
    localparam width_c3_conv_layer2_b                              = 64;
    localparam width_c3_conv_layer2_db                             = 64;
    localparam width_c3_conv_layer2_W                              = 64;
    localparam width_c3_conv_layer2_dW                             = 64;
    localparam width_c3_conv_layer2_map_common                     = 64;
    //struct:localparam width_s4_pooling_layer2                             = 21953536;
    localparam width_s4_pooling_layer2_data                        = 64;
    localparam width_s4_pooling_layer2_error                       = 64;
    localparam width_s4_pooling_layer2_b                           = 64;
    localparam width_s4_pooling_layer2_db                          = 64;
    localparam width_s4_pooling_layer2_W                           = 64;
    localparam width_s4_pooling_layer2_dW                          = 64;
    localparam width_s4_pooling_layer2_map_common                  = 64;
    //struct:localparam width_c5_conv_layer2                                = 21953536;
    localparam width_c5_conv_layer2_data                           = 64;
    localparam width_c5_conv_layer2_error                          = 64;
    localparam width_c5_conv_layer2_b                              = 64;
    localparam width_c5_conv_layer2_db                             = 64;
    localparam width_c5_conv_layer2_W                              = 64;
    localparam width_c5_conv_layer2_dW                             = 64;
    localparam width_c5_conv_layer2_map_common                     = 64;
    //struct:localparam width_output_layer2                                 = 21953536;
    localparam width_output_layer2_data                            = 64;
    localparam width_output_layer2_error                           = 64;
    localparam width_output_layer2_b                               = 64;
    localparam width_output_layer2_db                              = 64;
    localparam width_output_layer2_W                               = 64;
    localparam width_output_layer2_dW                              = 64;
    localparam width_output_layer2_map_common                      = 64;
    localparam width_pconnection                                   = 8;
    localparam width_generic_xmem32                                = 32;

    //xmem offset
    //struct:localparam offset_input_layer1                                 = 0;
    localparam offset_input_layer1_map_w                           = 0;
    localparam offset_input_layer1_map_h                           = 4;
    localparam offset_input_layer1_map_count                       = 8;
    localparam offset_input_layer1_kernel_w                        = 12;
    localparam offset_input_layer1_kernel_h                        = 16;
    localparam offset_input_layer1_kernel_count                    = 20;
    //struct:localparam offset_c1_conv_layer1                               = 24;
    localparam offset_c1_conv_layer1_map_w                         = 24;
    localparam offset_c1_conv_layer1_map_h                         = 28;
    localparam offset_c1_conv_layer1_map_count                     = 32;
    localparam offset_c1_conv_layer1_kernel_w                      = 36;
    localparam offset_c1_conv_layer1_kernel_h                      = 40;
    localparam offset_c1_conv_layer1_kernel_count                  = 44;
    //struct:localparam offset_s2_pooling_layer1                            = 48;
    localparam offset_s2_pooling_layer1_map_w                      = 48;
    localparam offset_s2_pooling_layer1_map_h                      = 52;
    localparam offset_s2_pooling_layer1_map_count                  = 56;
    localparam offset_s2_pooling_layer1_kernel_w                   = 60;
    localparam offset_s2_pooling_layer1_kernel_h                   = 64;
    localparam offset_s2_pooling_layer1_kernel_count               = 68;
    //struct:localparam offset_c3_conv_layer1                               = 72;
    localparam offset_c3_conv_layer1_map_w                         = 72;
    localparam offset_c3_conv_layer1_map_h                         = 76;
    localparam offset_c3_conv_layer1_map_count                     = 80;
    localparam offset_c3_conv_layer1_kernel_w                      = 84;
    localparam offset_c3_conv_layer1_kernel_h                      = 88;
    localparam offset_c3_conv_layer1_kernel_count                  = 92;
    //struct:localparam offset_s4_pooling_layer1                            = 96;
    localparam offset_s4_pooling_layer1_map_w                      = 96;
    localparam offset_s4_pooling_layer1_map_h                      = 100;
    localparam offset_s4_pooling_layer1_map_count                  = 104;
    localparam offset_s4_pooling_layer1_kernel_w                   = 108;
    localparam offset_s4_pooling_layer1_kernel_h                   = 112;
    localparam offset_s4_pooling_layer1_kernel_count               = 116;
    //struct:localparam offset_c5_conv_layer1                               = 120;
    localparam offset_c5_conv_layer1_map_w                         = 120;
    localparam offset_c5_conv_layer1_map_h                         = 124;
    localparam offset_c5_conv_layer1_map_count                     = 128;
    localparam offset_c5_conv_layer1_kernel_w                      = 132;
    localparam offset_c5_conv_layer1_kernel_h                      = 136;
    localparam offset_c5_conv_layer1_kernel_count                  = 140;
    //struct:localparam offset_output_layer1                                = 144;
    localparam offset_output_layer1_map_w                          = 144;
    localparam offset_output_layer1_map_h                          = 148;
    localparam offset_output_layer1_map_count                      = 152;
    localparam offset_output_layer1_kernel_w                       = 156;
    localparam offset_output_layer1_kernel_h                       = 160;
    localparam offset_output_layer1_kernel_count                   = 164;
    localparam offset_xxxxx_paddingA                               = 168;
    //struct:localparam offset_input_layer2                                 = 2048;
    localparam offset_input_layer2_data                            = 2048;
    localparam offset_input_layer2_error                           = 985088;
    localparam offset_input_layer2_b                               = 1968128;
    localparam offset_input_layer2_db                              = 1969088;
    localparam offset_input_layer2_W                               = 1970048;
    localparam offset_input_layer2_dW                              = 2354048;
    localparam offset_input_layer2_map_common                      = 2738048;
    //struct:localparam offset_c1_conv_layer2                               = 2746240;
    localparam offset_c1_conv_layer2_data                          = 2746240;
    localparam offset_c1_conv_layer2_error                         = 3729280;
    localparam offset_c1_conv_layer2_b                             = 4712320;
    localparam offset_c1_conv_layer2_db                            = 4713280;
    localparam offset_c1_conv_layer2_W                             = 4714240;
    localparam offset_c1_conv_layer2_dW                            = 5098240;
    localparam offset_c1_conv_layer2_map_common                    = 5482240;
    //struct:localparam offset_s2_pooling_layer2                            = 5490432;
    localparam offset_s2_pooling_layer2_data                       = 5490432;
    localparam offset_s2_pooling_layer2_error                      = 6473472;
    localparam offset_s2_pooling_layer2_b                          = 7456512;
    localparam offset_s2_pooling_layer2_db                         = 7457472;
    localparam offset_s2_pooling_layer2_W                          = 7458432;
    localparam offset_s2_pooling_layer2_dW                         = 7842432;
    localparam offset_s2_pooling_layer2_map_common                 = 8226432;
    //struct:localparam offset_c3_conv_layer2                               = 8234624;
    localparam offset_c3_conv_layer2_data                          = 8234624;
    localparam offset_c3_conv_layer2_error                         = 9217664;
    localparam offset_c3_conv_layer2_b                             = 10200704;
    localparam offset_c3_conv_layer2_db                            = 10201664;
    localparam offset_c3_conv_layer2_W                             = 10202624;
    localparam offset_c3_conv_layer2_dW                            = 10586624;
    localparam offset_c3_conv_layer2_map_common                    = 10970624;
    //struct:localparam offset_s4_pooling_layer2                            = 10978816;
    localparam offset_s4_pooling_layer2_data                       = 10978816;
    localparam offset_s4_pooling_layer2_error                      = 11961856;
    localparam offset_s4_pooling_layer2_b                          = 12944896;
    localparam offset_s4_pooling_layer2_db                         = 12945856;
    localparam offset_s4_pooling_layer2_W                          = 12946816;
    localparam offset_s4_pooling_layer2_dW                         = 13330816;
    localparam offset_s4_pooling_layer2_map_common                 = 13714816;
    //struct:localparam offset_c5_conv_layer2                               = 13723008;
    localparam offset_c5_conv_layer2_data                          = 13723008;
    localparam offset_c5_conv_layer2_error                         = 14706048;
    localparam offset_c5_conv_layer2_b                             = 15689088;
    localparam offset_c5_conv_layer2_db                            = 15690048;
    localparam offset_c5_conv_layer2_W                             = 15691008;
    localparam offset_c5_conv_layer2_dW                            = 16075008;
    localparam offset_c5_conv_layer2_map_common                    = 16459008;
    //struct:localparam offset_output_layer2                                = 16467200;
    localparam offset_output_layer2_data                           = 16467200;
    localparam offset_output_layer2_error                          = 17450240;
    localparam offset_output_layer2_b                              = 18433280;
    localparam offset_output_layer2_db                             = 18434240;
    localparam offset_output_layer2_W                              = 18435200;
    localparam offset_output_layer2_dW                             = 18819200;
    localparam offset_output_layer2_map_common                     = 19203200;
    localparam offset_pconnection                                  = 19211392;
    localparam offset_generic_xmem32                               = 0;

    //xmem depth
    //struct:localparam depth_input_layer1                                  = 1;
    localparam depth_input_layer1_map_w                            = 1;
    localparam depth_input_layer1_map_h                            = 1;
    localparam depth_input_layer1_map_count                        = 1;
    localparam depth_input_layer1_kernel_w                         = 1;
    localparam depth_input_layer1_kernel_h                         = 1;
    localparam depth_input_layer1_kernel_count                     = 1;
    //struct:localparam depth_c1_conv_layer1                                = 1;
    localparam depth_c1_conv_layer1_map_w                          = 1;
    localparam depth_c1_conv_layer1_map_h                          = 1;
    localparam depth_c1_conv_layer1_map_count                      = 1;
    localparam depth_c1_conv_layer1_kernel_w                       = 1;
    localparam depth_c1_conv_layer1_kernel_h                       = 1;
    localparam depth_c1_conv_layer1_kernel_count                   = 1;
    //struct:localparam depth_s2_pooling_layer1                             = 1;
    localparam depth_s2_pooling_layer1_map_w                       = 1;
    localparam depth_s2_pooling_layer1_map_h                       = 1;
    localparam depth_s2_pooling_layer1_map_count                   = 1;
    localparam depth_s2_pooling_layer1_kernel_w                    = 1;
    localparam depth_s2_pooling_layer1_kernel_h                    = 1;
    localparam depth_s2_pooling_layer1_kernel_count                = 1;
    //struct:localparam depth_c3_conv_layer1                                = 1;
    localparam depth_c3_conv_layer1_map_w                          = 1;
    localparam depth_c3_conv_layer1_map_h                          = 1;
    localparam depth_c3_conv_layer1_map_count                      = 1;
    localparam depth_c3_conv_layer1_kernel_w                       = 1;
    localparam depth_c3_conv_layer1_kernel_h                       = 1;
    localparam depth_c3_conv_layer1_kernel_count                   = 1;
    //struct:localparam depth_s4_pooling_layer1                             = 1;
    localparam depth_s4_pooling_layer1_map_w                       = 1;
    localparam depth_s4_pooling_layer1_map_h                       = 1;
    localparam depth_s4_pooling_layer1_map_count                   = 1;
    localparam depth_s4_pooling_layer1_kernel_w                    = 1;
    localparam depth_s4_pooling_layer1_kernel_h                    = 1;
    localparam depth_s4_pooling_layer1_kernel_count                = 1;
    //struct:localparam depth_c5_conv_layer1                                = 1;
    localparam depth_c5_conv_layer1_map_w                          = 1;
    localparam depth_c5_conv_layer1_map_h                          = 1;
    localparam depth_c5_conv_layer1_map_count                      = 1;
    localparam depth_c5_conv_layer1_kernel_w                       = 1;
    localparam depth_c5_conv_layer1_kernel_h                       = 1;
    localparam depth_c5_conv_layer1_kernel_count                   = 1;
    //struct:localparam depth_output_layer1                                 = 1;
    localparam depth_output_layer1_map_w                           = 1;
    localparam depth_output_layer1_map_h                           = 1;
    localparam depth_output_layer1_map_count                       = 1;
    localparam depth_output_layer1_kernel_w                        = 1;
    localparam depth_output_layer1_kernel_h                        = 1;
    localparam depth_output_layer1_kernel_count                    = 1;
    localparam depth_xxxxx_paddingA                                = 1880;
    //struct:localparam depth_input_layer2                                  = 1;
    localparam depth_input_layer2_data                             = 122880;
    localparam depth_input_layer2_error                            = 122880;
    localparam depth_input_layer2_b                                = 120;
    localparam depth_input_layer2_db                               = 120;
    localparam depth_input_layer2_W                                = 48000;
    localparam depth_input_layer2_dW                               = 48000;
    localparam depth_input_layer2_map_common                       = 1024;
    //struct:localparam depth_c1_conv_layer2                                = 1;
    localparam depth_c1_conv_layer2_data                           = 122880;
    localparam depth_c1_conv_layer2_error                          = 122880;
    localparam depth_c1_conv_layer2_b                              = 120;
    localparam depth_c1_conv_layer2_db                             = 120;
    localparam depth_c1_conv_layer2_W                              = 48000;
    localparam depth_c1_conv_layer2_dW                             = 48000;
    localparam depth_c1_conv_layer2_map_common                     = 1024;
    //struct:localparam depth_s2_pooling_layer2                             = 1;
    localparam depth_s2_pooling_layer2_data                        = 122880;
    localparam depth_s2_pooling_layer2_error                       = 122880;
    localparam depth_s2_pooling_layer2_b                           = 120;
    localparam depth_s2_pooling_layer2_db                          = 120;
    localparam depth_s2_pooling_layer2_W                           = 48000;
    localparam depth_s2_pooling_layer2_dW                          = 48000;
    localparam depth_s2_pooling_layer2_map_common                  = 1024;
    //struct:localparam depth_c3_conv_layer2                                = 1;
    localparam depth_c3_conv_layer2_data                           = 122880;
    localparam depth_c3_conv_layer2_error                          = 122880;
    localparam depth_c3_conv_layer2_b                              = 120;
    localparam depth_c3_conv_layer2_db                             = 120;
    localparam depth_c3_conv_layer2_W                              = 48000;
    localparam depth_c3_conv_layer2_dW                             = 48000;
    localparam depth_c3_conv_layer2_map_common                     = 1024;
    //struct:localparam depth_s4_pooling_layer2                             = 1;
    localparam depth_s4_pooling_layer2_data                        = 122880;
    localparam depth_s4_pooling_layer2_error                       = 122880;
    localparam depth_s4_pooling_layer2_b                           = 120;
    localparam depth_s4_pooling_layer2_db                          = 120;
    localparam depth_s4_pooling_layer2_W                           = 48000;
    localparam depth_s4_pooling_layer2_dW                          = 48000;
    localparam depth_s4_pooling_layer2_map_common                  = 1024;
    //struct:localparam depth_c5_conv_layer2                                = 1;
    localparam depth_c5_conv_layer2_data                           = 122880;
    localparam depth_c5_conv_layer2_error                          = 122880;
    localparam depth_c5_conv_layer2_b                              = 120;
    localparam depth_c5_conv_layer2_db                             = 120;
    localparam depth_c5_conv_layer2_W                              = 48000;
    localparam depth_c5_conv_layer2_dW                             = 48000;
    localparam depth_c5_conv_layer2_map_common                     = 1024;
    //struct:localparam depth_output_layer2                                 = 1;
    localparam depth_output_layer2_data                            = 122880;
    localparam depth_output_layer2_error                           = 122880;
    localparam depth_output_layer2_b                               = 120;
    localparam depth_output_layer2_db                              = 120;
    localparam depth_output_layer2_W                               = 48000;
    localparam depth_output_layer2_dW                              = 48000;
    localparam depth_output_layer2_map_common                      = 1024;
    localparam depth_pconnection                                   = 96;
    localparam depth_generic_xmem32                                = 4802872;

endpackage
